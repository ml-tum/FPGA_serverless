hyperloglog_wrapper hll_wrapper_inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .axi_ctrl(axi_ctrl),
    .axis_host_0_sink(axis_host_0_sink),
    .axis_host_0_src(axis_host_0_src)
    );
